module stats(
    input wire clk, // 27 MHz clock
    input wire reset, // reset
    input wire [7:0] inputs,
    input wire [4:0] random,
    output reg [3:0] hunger,
    output reg [3:0] happiness,
    output reg [3:0] health,
    output reg [3:0] hygiene,
    output reg [3:0] energy,
    // output reg [3:0] social
);

reg [26:0] count = 0;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        // Initialize all stats including social to 0 on reset
        hunger <= 4'd0;
        happiness <= 4'd0;
        health <= 4'd0;
        hygiene <= 4'd0;
        energy <= 4'd0;
        //social <= 4'd0;
    end else begin
        if (count == 27'd10_000_000) begin
            count <= 0;
            case (random)
                5'd0: begin
                    if (hunger < 4'd15) begin
                        hunger <= hunger + 1;
                    end
                end
                5'd1: begin
                    if (happiness < 4'd15) begin
                        happiness <= happiness + 1;
                    end
                end
                5'd2: begin
                    if (health < 4'd15) begin
                        health <= health + 1;
                    end
                end
                5'd3: begin
                    if (hygiene < 4'd15) begin
                        hygiene <= hygiene + 1;
                    end
                end
                5'd4: begin
                    if (energy < 4'd15) begin
                        energy <= energy + 1;
                    end
                end
                // 5'd5: begin
                //     if (social < 4'd15) begin
                //         social <= social + 1;
                //     end
                // end
            endcase
        end
        else begin
            count <= count + 1;
        end
    end
end

// logic to decrease stats
always @(posedge clk or posedge reset) begin
    if (reset) begin
        // Reset the stats to 0 on reset
        hunger <= 4'd0;
        happiness <= 4'd0;
        health <= 4'd0;
        hygiene <= 4'd0;
        energy <= 4'd0;
        // social <= 4'd0;
    end else begin
        if (inputs[0] == 1'b1) begin
            if (hunger > 4'd0) begin
                hunger <= hunger - 1;
            end
        end
        if (inputs[1] == 1'b1) begin
            if (happiness > 4'd0) begin
                happiness <= happiness - 1;
            end
        end
        if (inputs[2] == 1'b1) begin
            if (health > 4'd0) begin
                health <= health - 1;
            end
        end
        if (inputs[3] == 1'b1) begin
            if (hygiene > 4'd0) begin
                hygiene <= hygiene - 1;
            end
        end
        if (inputs[4] == 1'b1) begin
            if (energy > 4'd0) begin
                energy <= energy - 1;
            end
        end
        // if (inputs[5] == 1'b1) begin
        //     if (social > 4'd0) begin
        //         social <= social - 1;
        //     end
        // end
    end
end

endmodule
